`define ARTY_A7

`define ARIANE_DATA_WIDTH 64

// Instantiate protocl checker
// `define PROTOCOL_CHECKER

// write-back cache
// `define WB_DCACHE

// write-through cache
`define WT_DCACHE

`define RAMB16

// include NEXYS_VIDEO specific code (DDR3, clock gen, leds/sw)
// `define NEXYS_VIDEO